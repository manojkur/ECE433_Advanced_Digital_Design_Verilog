module ControlUnit (
	input clock,
	input ClockI2C,
	input Go,
	input Reset,
	output BaudEnable,
	output ReadorWrite,
	ouptut Select,
	output ShiftorHold,
	output StartStopAck,
	output WriteLoad,	
);




endmodule