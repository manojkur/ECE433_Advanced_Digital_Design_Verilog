module I2C__SDAmodule (
	inout SDA,
	input ReadOrWrite,
	input Select,
	input StartStopAck,
	output ShiftDataIn,
	input ShiftDataOut));



endmodule