module I2C_SDAmodule (
	inout SDA,
	input ReadOrWrite,
	input Select,
	input StartStopAck,
	output ShiftDataIn,
	input ShiftDataOut);



endmodule